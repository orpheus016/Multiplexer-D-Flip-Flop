* Inverter Testbench

* Include the sky130 model library
.lib "/foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice" tt

* Include the extracted netlist for the inverter
.include "/foss/designs/UTS/Gates/Inverter/inverter.spice"

* Sumber Tegangan (Voltage Sources)
Vpwr Vpwr 0 DC 1.8
Vgnd Vgnd 0 DC 0

* Input Pulse Source
VIN IN 0 PULSE(0 1.8 0 10p 10p 10n 20n)

* Inverter Instantiation
Xinv IN OUT Vpwr Vgnd Inverter

* Perintah Simulasi Transien
.tran 0.1n 40n

* Perintah untuk Output
.control
  run
  plot v(IN)+2 v(OUT)
.endc

.end

