magic
tech sky130A
timestamp 1745050697
<< error_s >>
rect 296 330 305 370
rect 310 330 319 370
<< nwell >>
rect 895 375 905 715
<< metal1 >>
rect 0 695 905 725
rect 65 330 305 370
rect 310 330 345 370
rect 415 330 480 370
rect 720 295 760 330
rect 145 255 185 295
rect 240 270 245 295
rect 210 240 245 270
rect 560 255 600 295
rect 655 255 760 295
rect 865 255 900 295
rect 210 210 215 240
rect 210 205 245 210
rect 800 240 840 255
rect 800 210 805 240
rect 835 210 840 240
rect 800 205 840 210
rect 0 0 905 30
<< via1 >>
rect 215 210 245 240
rect 805 210 835 240
<< metal2 >>
rect 210 240 840 245
rect 210 210 215 240
rect 245 210 805 240
rect 835 210 840 240
rect 210 205 840 210
use inverter  inverter_0
timestamp 1744986694
transform 1 0 345 0 1 195
box -105 -195 80 530
use nand  nand_0
timestamp 1744987844
transform 1 0 105 0 1 195
box -105 -195 145 530
use nand  nand_1
timestamp 1744987844
transform 1 0 520 0 1 195
box -105 -195 145 530
use nand  nand_2
timestamp 1744987844
transform 1 0 760 0 1 195
box -105 -195 145 530
<< labels >>
flabel metal1 865 255 900 295 1 FreeSans 200 0 0 0 D
port 6 n
flabel metal1 0 0 905 30 1 FreeSans 200 0 0 0 Vgnd
port 5 n
flabel metal1 0 695 905 725 1 FreeSans 200 0 0 0 Vpwr
port 4 n
flabel metal1 75 340 95 360 1 FreeSans 200 0 0 0 S
port 1 n
flabel metal1 560 255 600 295 1 FreeSans 200 0 0 0 A
port 2 n
flabel metal1 145 255 185 295 1 FreeSans 200 0 0 0 B
port 3 n
<< end >>
