magic
tech sky130A
timestamp 1744986694
<< nwell >>
rect -105 180 80 520
<< nmos >>
rect 0 -150 15 50
<< pmos >>
rect 0 200 15 500
<< ndiff >>
rect -45 35 0 50
rect -45 -35 -35 35
rect -15 -35 0 35
rect -45 -65 0 -35
rect -45 -135 -35 -65
rect -15 -135 0 -65
rect -45 -150 0 -135
rect 15 35 60 50
rect 15 -35 30 35
rect 50 -35 60 35
rect 15 -65 60 -35
rect 15 -135 30 -65
rect 50 -135 60 -65
rect 15 -150 60 -135
<< pdiff >>
rect -45 485 0 500
rect -45 415 -35 485
rect -15 415 0 485
rect -45 385 0 415
rect -45 315 -35 385
rect -15 315 0 385
rect -45 285 0 315
rect -45 215 -35 285
rect -15 215 0 285
rect -45 200 0 215
rect 15 485 60 500
rect 15 415 30 485
rect 50 415 60 485
rect 15 385 60 415
rect 15 315 30 385
rect 50 315 60 385
rect 15 285 60 315
rect 15 215 30 285
rect 50 215 60 285
rect 15 200 60 215
<< ndiffc >>
rect -35 -35 -15 35
rect -35 -135 -15 -65
rect 30 -35 50 35
rect 30 -135 50 -65
<< pdiffc >>
rect -35 415 -15 485
rect -35 315 -15 385
rect -35 215 -15 285
rect 30 415 50 485
rect 30 315 50 385
rect 30 215 50 285
<< psubdiff >>
rect -85 35 -45 50
rect -85 -35 -75 35
rect -55 -35 -45 35
rect -85 -65 -45 -35
rect -85 -135 -75 -65
rect -55 -135 -45 -65
rect -85 -150 -45 -135
<< nsubdiff >>
rect -85 485 -45 500
rect -85 415 -75 485
rect -55 415 -45 485
rect -85 385 -45 415
rect -85 315 -75 385
rect -55 315 -45 385
rect -85 285 -45 315
rect -85 215 -75 285
rect -55 215 -45 285
rect -85 200 -45 215
<< psubdiffcont >>
rect -75 -35 -55 35
rect -75 -135 -55 -65
<< nsubdiffcont >>
rect -75 415 -55 485
rect -75 315 -55 385
rect -75 215 -55 285
<< poly >>
rect 0 500 15 515
rect 0 100 15 200
rect -40 90 15 100
rect -40 70 -30 90
rect -10 70 15 90
rect -40 60 15 70
rect 0 50 15 60
rect 0 -165 15 -150
<< polycont >>
rect -30 70 -10 90
<< locali >>
rect -85 525 -65 530
rect -85 490 -65 505
rect -85 485 -5 490
rect -85 415 -75 485
rect -55 415 -35 485
rect -15 415 -5 485
rect -85 410 -5 415
rect 20 485 60 490
rect 20 415 30 485
rect 50 415 60 485
rect 20 410 60 415
rect -85 390 -65 410
rect 40 390 60 410
rect -85 385 -5 390
rect -85 315 -75 385
rect -55 315 -35 385
rect -15 315 -5 385
rect -85 310 -5 315
rect 20 385 60 390
rect 20 315 30 385
rect 50 315 60 385
rect 20 310 60 315
rect -85 290 -65 310
rect 40 290 60 310
rect -85 285 -5 290
rect -85 215 -75 285
rect -55 215 -35 285
rect -15 215 -5 285
rect -85 210 -5 215
rect 20 285 60 290
rect 20 215 30 285
rect 50 215 60 285
rect 20 210 60 215
rect -40 90 0 100
rect -40 70 -30 90
rect -10 70 0 90
rect -40 60 0 70
rect 40 95 60 210
rect 40 90 65 95
rect 40 70 45 90
rect 40 65 65 70
rect 40 40 60 65
rect -85 35 -5 40
rect -85 -35 -75 35
rect -55 -35 -35 35
rect -15 -35 -5 35
rect -85 -40 -5 -35
rect 20 35 60 40
rect 20 -35 30 35
rect 50 -35 60 35
rect 20 -40 60 -35
rect -85 -60 -65 -40
rect 40 -60 60 -40
rect -85 -65 -5 -60
rect -85 -135 -75 -65
rect -55 -135 -35 -65
rect -15 -135 -5 -65
rect -85 -140 -5 -135
rect 20 -65 60 -60
rect 20 -135 30 -65
rect 50 -135 60 -65
rect 20 -140 60 -135
rect -85 -170 -65 -140
rect -85 -195 -65 -190
<< viali >>
rect -85 505 -65 525
rect -30 70 -10 90
rect 45 70 65 90
rect -85 -190 -65 -170
<< metal1 >>
rect -105 525 80 530
rect -105 505 -85 525
rect -65 505 80 525
rect -105 500 80 505
rect -40 90 0 100
rect -40 70 -30 90
rect -10 70 0 90
rect -40 60 0 70
rect 40 90 75 100
rect 40 70 45 90
rect 65 70 75 90
rect 40 60 75 70
rect -105 -170 80 -165
rect -105 -190 -85 -170
rect -65 -190 80 -170
rect -105 -195 80 -190
<< labels >>
flabel viali -85 -190 -65 -170 1 FreeSans 200 0 0 0 Vgnd
port 4 n
flabel metal1 -30 70 -10 90 1 FreeSans 200 0 0 0 IN
port 1 n
flabel viali -85 505 -65 525 1 FreeSans 200 0 0 0 Vpwr
port 3 n
flabel metal1 40 60 75 100 1 FreeSans 200 0 0 0 OUT
port 2 n
<< end >>
