* Inverter Testbench

* Include the sky130 model library
.lib "/foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice" tt

* Include the extracted netlist for the inverter
.include "/foss/designs/UTS/Gates/NAND/nand.spice"

* Sumber Tegangan (Voltage Sources)
Vpwr Vpwr 0 DC 1.8
Vgnd Vgnd 0 DC 0

* Input Pulse Source
VINA A 0 PULSE(0 1.8 0 10p 10p 10n 20n)
VINB B 0 PULSE(0 1.8 0 10p 10p 20n 40n)

* Inverter Instantiation
Xnand A OUT Vpwr Vgnd B nand

* Perintah Simulasi Transien
.tran 0.1n 40n

* Perintah untuk Output
.control
  run
  plot v(A)+4 v(B)+2 v(OUT)
.endc

.end

